LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LAB305 IS
	PORT(SW: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		  HEX0: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		  HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		  HEX2: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		  HEX3: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		  KEY: IN STD_LOGIC_VECTOR(2 DOWNTO 0));
END LAB305;

ARCHITECTURE Behavior OF LAB305 IS 
	COMPONENT char_7seg
		PORT ( V : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				 Display : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
	END COMPONENT;

SIGNAL Resetn: STD_LOGIC;
SIGNAL CLK: STD_LOGIC;
SIGNAL D: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL Q: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL S: STD_LOGIC;
SIGNAL A: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL B: STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN 

	Resetn <= KEY(0);
	CLK <= KEY(1);
	D <= SW(7 DOWNTO 0);
	S <= SW(9);

	PROCESS(Resetn, CLK, SW)
	BEGIN 
		IF Resetn = '0' THEN
			Q <= "00000000";
		ELSIF CLK'EVENT AND CLK = '1' THEN
			Q <= D;
		END IF;
	END PROCESS;
	
	PROCESS(S, Q)
	BEGIN 
		IF S = '0' THEN
			A <= Q;
		ELSIF S = '1' THEN
			B <= Q;
		END IF;
	END PROCESS;
	
	
	
	M0:char_7seg PORT MAP (A(3 DOWNTO 0), HEX2);
	M1:char_7seg PORT MAP (A(7 DOWNTO 4), HEX3);
		
	M2:char_7seg PORT MAP (B(3 DOWNTO 0), HEX0);
	M3:char_7seg PORT MAP (B(7 DOWNTO 4), HEX1);
	

END Behavior;



LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY char_7seg IS
	PORT ( V : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 Display : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END char_7seg;

ARCHITECTURE Behavior OF char_7seg IS
BEGIN
	WITH V SELECT
		Display <= "1000000" WHEN "0000",--0
					  "1111001" WHEN "0001",--1
						"0100100" WHEN "0010",--2
						"0110000" WHEN "0011",--3
						"0011001" WHEN "0100",--4
						"0010010" WHEN "0101",--5
						"0000010" WHEN "0110",--6
						"1011000" WHEN "0111",--7
						"0000000" WHEN "1000",--8
						"0010000" WHEN "1001",--9
						"0001000" WHEN "1010",--A
						"0000011" WHEN "1011",--b
						"1000110" WHEN "1100",--C
						"0100001" WHEN "1101",--d
						"0000110" WHEN "1110",--E
						"0001110" WHEN "1111";--F
END Behavior;



