library verilog;
use verilog.vl_types.all;
entity LAB901_vlg_vec_tst is
end LAB901_vlg_vec_tst;
