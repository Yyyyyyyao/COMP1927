library verilog;
use verilog.vl_types.all;
entity LAB501_vlg_vec_tst is
end LAB501_vlg_vec_tst;
