LIBRARY ieee; 
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;


ENTITY EX1 IS 
	PORT(A: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		  B: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		  RESULT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END EX1;

ARCHITECTURE Behavior OF EX1 IS

SIGNAL P: STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL Q: STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL SUB: STD_LOGIC_VECTOR(10 DOWNTO 0);

BEGIN 

	P <= '0' & A;
	Q <= '0' & B;
	
	SUB <= P + (NOT(Q) + '1');
	RESULT <= SUB(10 DOWNTO 8);


END Behavior; 
