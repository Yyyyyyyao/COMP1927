cmp16_inst : cmp16 PORT MAP (
		dataa	 => dataa_sig,
		alb	 => alb_sig
	);
