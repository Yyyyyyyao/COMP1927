LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LAB204 IS
PORT ( SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 HEX3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);		 
		 LEDR: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		 LEDG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END LAB204;

ARCHITECTURE Behavior OF LAB204 IS
	COMPONENT comparator
	PORT ( U : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 Cout: IN STD_LOGIC;
			 z : OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT char_7seg
		PORT ( C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				Display0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT circuit_a
		PORT ( A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				 B: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT mul_2to1
		PORT ( B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				 V : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				 s : IN STD_LOGIC;
				 M: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT circuit_b
			PORT (s : IN STD_LOGIC;
					K: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT full_adder
		PORT (Cin, x, y: IN STD_LOGIC;
				s, Cout: OUT STD_LOGIC);
	END COMPONENT;
	
	
SIGNAL M : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL V : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL O : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL z : STD_LOGIC;


SIGNAL C: STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL A: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL B: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL S: STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	
	
BEGIN
	
	LEDR <= SW;
	C(0) <= SW(8);
	A <= SW(7 DOWNTO 4);
	B <= SW(3 DOWNTO 0);
	LEDG(4) <= C(4);
	LEDG(0) <= S(0); 
	LEDG(1) <= S(1); 
	LEDG(2) <= S(2);
	LEDG(3) <= S(3);
	
	
	step0: full_adder PORT MAP(C(0), A(0), B(0), S(0), C(1));
	step1: full_adder PORT MAP(C(1), A(1), B(1), S(1), C(2));
	step2: full_adder PORT MAP(C(2), A(2), B(2), S(2), C(3));
	step3: full_adder PORT MAP(C(3), A(3), B(3), S(3), C(4));
	
	V <= S;
	M0: comparator PORT MAP (V, C(4),z);
	M1: circuit_a PORT MAP (V, O);
	M2: mul_2to1 PORT MAP (O, V, z, M);
	M3: char_7seg PORT MAP (M, HEX0);
	M4: circuit_b PORT MAP (z, HEX1);
	M5: char_7seg PORT MAP (A, HEX3);
	M6: char_7seg PORT MAP (B, HEX2);
	
	LEDG(7) <= (A(1) AND A(3)) OR (A(2) AND A(3)) OR (B(1) AND B(3)) OR (B(2) AND B(3));
	
END Behavior;

--full_adder
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY full_adder IS
	PORT (Cin, x, y: IN STD_LOGIC;
			s, Cout: OUT STD_LOGIC);
END full_adder;

ARCHITECTURE Behavior OF full_adder IS
BEGIN
	s <= x XOR y XOR Cin;
	Cout <= (x AND y) OR (Cin AND x) OR (Cin AND y);


END Behavior;

--Circuit_B
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY circuit_b IS
	PORT (s: IN STD_LOGIC;
			K: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END circuit_b;

ARCHITECTURE Behavior OF circuit_b IS
BEGIN
	K(0) <= s;
	K(1) <= '0';
	K(2) <= '0';
	K(3) <= s;
	K(4) <= s;
	K(5) <= s;
	K(6) <= '1';


END Behavior;




--mul_2to1
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mul_2to1 IS
	PORT ( B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 V : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 s : IN STD_LOGIC;
			 M: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END mul_2to1;

ARCHITECTURE Behavior OF mul_2to1 IS
BEGIN

	M(0) <= (s AND B(0)) OR (NOT(s) AND V(0));
	M(1) <= (s AND B(1)) OR (NOT(s) AND V(1));
	M(2) <= (s AND B(2)) OR (NOT(s) AND V(2));
	M(3) <= (s AND B(3)) OR (NOT(s) AND V(3));
	
END Behavior;





--Circuit_A
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY circuit_a IS
	PORT ( A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 B: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END circuit_a;

ARCHITECTURE Behavior OF circuit_a IS
BEGIN
	B(3) <= A(1) AND NOT(A(3)) AND NOT(A(2));
	B(2) <= (A(1) AND A(2) AND A(3)) OR (NOT A(1) AND NOT A(2) AND NOT A(3));
	B(1) <= NOT(A(1));
	B(0) <= A(0);
END Behavior;



--Comparator
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY comparator IS
	PORT ( U : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 Cout: IN STD_LOGIC;
			 z : OUT STD_LOGIC);
END comparator;

ARCHITECTURE Behavior OF comparator IS
BEGIN
	z <= (U(2) AND U(3)) OR (U(1) AND U(3)) OR Cout;
	
END Behavior;




--7 segment decoder
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY char_7seg IS
	PORT ( C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 Display0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END char_7seg;

ARCHITECTURE Behavior OF char_7seg IS
BEGIN
	Display0(0) <= NOT(C(3) OR C(1) OR (C(2) AND C(0)) OR (NOT(C(2)) AND NOT(C(0))));
	Display0(1) <= NOT(NOT(C(2)) OR (NOT(C(1)) AND NOT(C(0))) OR (C(1) AND C(0)));
	Display0(2) <= NOT(C(2) OR NOT(C(1)) OR C(0));
	Display0(3) <= NOT((NOT(C(2)) AND NOT(C(0))) OR (C(1) AND NOT(C(0))) OR (C(2) AND NOT(C(1)) AND C(0)) OR (NOT(C(2)) AND C(1)) OR C(3));
	Display0(4) <= NOT((NOT(C(2)) AND NOT(C(0))) OR (C(1) AND NOT(C(0))));
	Display0(5) <= NOT(C(3) OR (NOT(C(1)) AND NOT(C(0))) OR (C(2) AND NOT(C(1))) OR (C(2) AND NOT(C(0))));
	Display0(6) <= NOT(C(3) OR (C(2) AND NOT(C(1))) OR (C(1) AND NOT(C(2))) OR (C(1) AND NOT(C(0))));
	
END Behavior;