compare_inst : compare PORT MAP (
		dataa	 => dataa_sig,
		agb	 => agb_sig
	);
