library verilog;
use verilog.vl_types.all;
entity LAB304_vlg_vec_tst is
end LAB304_vlg_vec_tst;
