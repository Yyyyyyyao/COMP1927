library verilog;
use verilog.vl_types.all;
entity LAB204_vlg_vec_tst is
end LAB204_vlg_vec_tst;
