compare11_inst : compare11 PORT MAP (
		dataa	 => dataa_sig,
		aeb	 => aeb_sig
	);
