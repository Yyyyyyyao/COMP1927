LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LAB302 IS

PORT ( Clk,D: IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END LAB302;

ARCHITECTURE Structural OF LAB302 IS

SIGNAL R_g, S_g, Qa, Qb : STD_LOGIC ;

ATTRIBUTE keep : boolean;
ATTRIBUTE keep of R_g, S_g, Qa, Qb : SIGNAL IS true;

BEGIN

S_g <= NOT(D AND Clk);
R_g <= NOT(NOT D AND Clk);
Qa <= NOT(S_g AND Qb);
Qb <= NOT(Qa AND R_g);


Q <= Qa;


END Structural;