compare16_inst : compare16 PORT MAP (
		dataa	 => dataa_sig,
		agb	 => agb_sig
	);
