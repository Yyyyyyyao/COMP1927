compare21_inst : compare21 PORT MAP (
		dataa	 => dataa_sig,
		agb	 => agb_sig
	);
