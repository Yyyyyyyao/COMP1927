library verilog;
use verilog.vl_types.all;
entity LAB401_vlg_vec_tst is
end LAB401_vlg_vec_tst;
