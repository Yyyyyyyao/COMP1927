LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LAB101 IS
	PORT ( SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
			LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END LAB101;

ARCHITECTURE Behavior OF LAB101 IS
BEGIN
	LEDR <= SW;
END Behavior;